`timescale 1ns / 1ps

module SectorProcessor(
  input clk,
  input reset,
  input en_proc,
  input[2:0] bx_in_MatchCalculator,
  output CM_L3PHIC20_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC20_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC20_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC20_nentries_0_V_dout,
  input[7:0] CM_L3PHIC20_nentries_1_V_dout,
  output CM_L3PHIC21_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC21_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC21_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC21_nentries_0_V_dout,
  input[7:0] CM_L3PHIC21_nentries_1_V_dout,
  output AS_L3PHICn4_dataarray_data_V_enb,
  output[9:0] AS_L3PHICn4_dataarray_data_V_readaddr,
  input[35:0] AS_L3PHICn4_dataarray_data_V_dout,
  input[7:0] AS_L3PHICn4_nentries_0_V_dout,
  input[7:0] AS_L3PHICn4_nentries_1_V_dout,
  input[7:0] AS_L3PHICn4_nentries_2_V_dout,
  input[7:0] AS_L3PHICn4_nentries_3_V_dout,
  input[7:0] AS_L3PHICn4_nentries_4_V_dout,
  input[7:0] AS_L3PHICn4_nentries_5_V_dout,
  input[7:0] AS_L3PHICn4_nentries_6_V_dout,
  input[7:0] AS_L3PHICn4_nentries_7_V_dout,
  output CM_L3PHIC22_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC22_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC22_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC22_nentries_0_V_dout,
  input[7:0] CM_L3PHIC22_nentries_1_V_dout,
  output CM_L3PHIC23_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC23_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC23_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC23_nentries_0_V_dout,
  input[7:0] CM_L3PHIC23_nentries_1_V_dout,
  output CM_L3PHIC24_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC24_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC24_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC24_nentries_0_V_dout,
  input[7:0] CM_L3PHIC24_nentries_1_V_dout,
  output CM_L3PHIC17_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC17_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC17_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC17_nentries_0_V_dout,
  input[7:0] CM_L3PHIC17_nentries_1_V_dout,
  output CM_L3PHIC18_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC18_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC18_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC18_nentries_0_V_dout,
  input[7:0] CM_L3PHIC18_nentries_1_V_dout,
  output AP_L3PHIC_dataarray_data_V_enb,
  output[9:0] AP_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] AP_L3PHIC_dataarray_data_V_dout,
  input[7:0] AP_L3PHIC_nentries_0_V_dout,
  input[7:0] AP_L3PHIC_nentries_1_V_dout,
  input[7:0] AP_L3PHIC_nentries_2_V_dout,
  input[7:0] AP_L3PHIC_nentries_3_V_dout,
  input[7:0] AP_L3PHIC_nentries_4_V_dout,
  input[7:0] AP_L3PHIC_nentries_5_V_dout,
  input[7:0] AP_L3PHIC_nentries_6_V_dout,
  input[7:0] AP_L3PHIC_nentries_7_V_dout,
  output CM_L3PHIC19_dataarray_data_V_enb,
  output[7:0] CM_L3PHIC19_dataarray_data_V_readaddr,
  input[13:0] CM_L3PHIC19_dataarray_data_V_dout,
  input[7:0] CM_L3PHIC19_nentries_0_V_dout,
  input[7:0] CM_L3PHIC19_nentries_1_V_dout,
  output[2:0] bx_out_MatchCalculator,
  output FM_L1L2XX_L3PHIC_dataarray_data_V_wea,
  output[7:0] FM_L1L2XX_L3PHIC_dataarray_data_V_writeaddr,
  output[44:0] FM_L1L2XX_L3PHIC_dataarray_data_V_din,
  output FM_L1L2XX_L3PHIC_nentries_0_V_we,
  output[7:0] FM_L1L2XX_L3PHIC_nentries_0_V_din,
  output FM_L1L2XX_L3PHIC_nentries_1_V_we,
  output[7:0] FM_L1L2XX_L3PHIC_nentries_1_V_din,
  output FM_L5L6XX_L3PHIC_dataarray_data_V_wea,
  output[7:0] FM_L5L6XX_L3PHIC_dataarray_data_V_writeaddr,
  output[44:0] FM_L5L6XX_L3PHIC_dataarray_data_V_din,
  output FM_L5L6XX_L3PHIC_nentries_0_V_we,
  output[7:0] FM_L5L6XX_L3PHIC_nentries_0_V_din,
  output FM_L5L6XX_L3PHIC_nentries_1_V_we,
  output[7:0] FM_L5L6XX_L3PHIC_nentries_1_V_din,
  output MatchCalculator_done
);

MatchCalculatorTop_0 MC_L3PHIC(
  .ap_clk(clk),
  .ap_rst(reset),
  .ap_start(en_proc),
  .ap_done(MatchCalculator_done),
  .bx_V(bx_in_MatchCalculator),
  .match1_dataarray_data_V_ce0(CM_L3PHIC17_dataarray_data_V_enb),
  .match1_dataarray_data_V_address0(CM_L3PHIC17_dataarray_data_V_readaddr),
  .match1_dataarray_data_V_q0(CM_L3PHIC17_dataarray_data_V_dout),
  .match1_nentries_0_V(CM_L3PHIC17_nentries_0_V_dout),
  .match1_nentries_1_V(CM_L3PHIC17_nentries_1_V_dout),
  .match2_dataarray_data_V_ce0(CM_L3PHIC18_dataarray_data_V_enb),
  .match2_dataarray_data_V_address0(CM_L3PHIC18_dataarray_data_V_readaddr),
  .match2_dataarray_data_V_q0(CM_L3PHIC18_dataarray_data_V_dout),
  .match2_nentries_0_V(CM_L3PHIC18_nentries_0_V_dout),
  .match2_nentries_1_V(CM_L3PHIC18_nentries_1_V_dout),
  .match3_dataarray_data_V_ce0(CM_L3PHIC19_dataarray_data_V_enb),
  .match3_dataarray_data_V_address0(CM_L3PHIC19_dataarray_data_V_readaddr),
  .match3_dataarray_data_V_q0(CM_L3PHIC19_dataarray_data_V_dout),
  .match3_nentries_0_V(CM_L3PHIC19_nentries_0_V_dout),
  .match3_nentries_1_V(CM_L3PHIC19_nentries_1_V_dout),
  .match4_dataarray_data_V_ce0(CM_L3PHIC20_dataarray_data_V_enb),
  .match4_dataarray_data_V_address0(CM_L3PHIC20_dataarray_data_V_readaddr),
  .match4_dataarray_data_V_q0(CM_L3PHIC20_dataarray_data_V_dout),
  .match4_nentries_0_V(CM_L3PHIC20_nentries_0_V_dout),
  .match4_nentries_1_V(CM_L3PHIC20_nentries_1_V_dout),
  .match5_dataarray_data_V_ce0(CM_L3PHIC21_dataarray_data_V_enb),
  .match5_dataarray_data_V_address0(CM_L3PHIC21_dataarray_data_V_readaddr),
  .match5_dataarray_data_V_q0(CM_L3PHIC21_dataarray_data_V_dout),
  .match5_nentries_0_V(CM_L3PHIC21_nentries_0_V_dout),
  .match5_nentries_1_V(CM_L3PHIC21_nentries_1_V_dout),
  .match6_dataarray_data_V_ce0(CM_L3PHIC22_dataarray_data_V_enb),
  .match6_dataarray_data_V_address0(CM_L3PHIC22_dataarray_data_V_readaddr),
  .match6_dataarray_data_V_q0(CM_L3PHIC22_dataarray_data_V_dout),
  .match6_nentries_0_V(CM_L3PHIC22_nentries_0_V_dout),
  .match6_nentries_1_V(CM_L3PHIC22_nentries_1_V_dout),
  .match7_dataarray_data_V_ce0(CM_L3PHIC23_dataarray_data_V_enb),
  .match7_dataarray_data_V_address0(CM_L3PHIC23_dataarray_data_V_readaddr),
  .match7_dataarray_data_V_q0(CM_L3PHIC23_dataarray_data_V_dout),
  .match7_nentries_0_V(CM_L3PHIC23_nentries_0_V_dout),
  .match7_nentries_1_V(CM_L3PHIC23_nentries_1_V_dout),
  .match8_dataarray_data_V_ce0(CM_L3PHIC24_dataarray_data_V_enb),
  .match8_dataarray_data_V_address0(CM_L3PHIC24_dataarray_data_V_readaddr),
  .match8_dataarray_data_V_q0(CM_L3PHIC24_dataarray_data_V_dout),
  .match8_nentries_0_V(CM_L3PHIC24_nentries_0_V_dout),
  .match8_nentries_1_V(CM_L3PHIC24_nentries_1_V_dout),
  .allstub_dataarray_data_V_ce0(AS_L3PHICn4_dataarray_data_V_enb),
  .allstub_dataarray_data_V_address0(AS_L3PHICn4_dataarray_data_V_readaddr),
  .allstub_dataarray_data_V_q0(AS_L3PHICn4_dataarray_data_V_dout),
  .allstub_nentries_V_q0(AS_L3PHICn4_nentries_0_V_dout),
  .allstub_nentries_V_q1(AS_L3PHICn4_nentries_1_V_dout),
  /*
  .allstub_nentries_V_q2(AS_L3PHICn4_nentries_2_V_dout),
  .allstub_nentries_V_q3(AS_L3PHICn4_nentries_3_V_dout),
  .allstub_nentries_V_q4(AS_L3PHICn4_nentries_4_V_dout),
  .allstub_nentries_V_q5(AS_L3PHICn4_nentries_5_V_dout),
  .allstub_nentries_V_q6(AS_L3PHICn4_nentries_6_V_dout),
  .allstub_nentries_V_q7(AS_L3PHICn4_nentries_7_V_dout),
  */
  .allproj_dataarray_data_V_ce0(AP_L3PHIC_dataarray_data_V_enb),
  .allproj_dataarray_data_V_address0(AP_L3PHIC_dataarray_data_V_readaddr),
  .allproj_dataarray_data_V_q0(AP_L3PHIC_dataarray_data_V_dout),
  .allproj_nentries_V_q0(AP_L3PHIC_nentries_0_V_dout),
  /*
  .allproj_nentries_V_q1(AP_L3PHIC_nentries_1_V_dout),
  .allproj_nentries_V_q2(AP_L3PHIC_nentries_2_V_dout),
  .allproj_nentries_V_q3(AP_L3PHIC_nentries_3_V_dout),
  .allproj_nentries_V_q4(AP_L3PHIC_nentries_4_V_dout),
  .allproj_nentries_V_q5(AP_L3PHIC_nentries_5_V_dout),
  .allproj_nentries_V_q6(AP_L3PHIC_nentries_6_V_dout),
  .allproj_nentries_V_q7(AP_L3PHIC_nentries_7_V_dout),
  */
  .bx_o_V(bx_out_MatchCalculator),
  .fullmatch1_dataarray_data_V_we0(FM_L1L2XX_L3PHIC_dataarray_data_V_wea),
  .fullmatch1_dataarray_data_V_address0(FM_L1L2XX_L3PHIC_dataarray_data_V_writeaddr),
  .fullmatch1_dataarray_data_V_d0(FM_L1L2XX_L3PHIC_dataarray_data_V_din),
  .fullmatch1_nentries_0_V_ap_vld(FM_L1L2XX_L3PHIC_nentries_0_V_we),
  .fullmatch1_nentries_0_V(FM_L1L2XX_L3PHIC_nentries_0_V_din),
  .fullmatch1_nentries_1_V_ap_vld(FM_L1L2XX_L3PHIC_nentries_1_V_we),
  .fullmatch1_nentries_1_V(FM_L1L2XX_L3PHIC_nentries_1_V_din),
  .fullmatch3_dataarray_data_V_we0(FM_L5L6XX_L3PHIC_dataarray_data_V_wea),
  .fullmatch3_dataarray_data_V_address0(FM_L5L6XX_L3PHIC_dataarray_data_V_writeaddr),
  .fullmatch3_dataarray_data_V_d0(FM_L5L6XX_L3PHIC_dataarray_data_V_din),
  .fullmatch3_nentries_0_V_ap_vld(FM_L5L6XX_L3PHIC_nentries_0_V_we),
  .fullmatch3_nentries_0_V(FM_L5L6XX_L3PHIC_nentries_0_V_din),
  .fullmatch3_nentries_1_V_ap_vld(FM_L5L6XX_L3PHIC_nentries_1_V_we),
  .fullmatch3_nentries_1_V(FM_L5L6XX_L3PHIC_nentries_1_V_din)
);

endmodule
